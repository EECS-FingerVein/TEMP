`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/09/2022 07:53:03 PM
// Design Name: 
// Module Name: reg_1C
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module reg_1C(addr, datain, dataout, sig);

    input [7:0] addr;
    input [8:0] datain;
    input sig;
    
    output [8:0] dataout;
    
    
    
endmodule
